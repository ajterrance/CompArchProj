module not_1b(x, o);
  
  output o;
  input x;
  
  assign o = !x;
  
endmodule
